`define INWVAL 24
`define RVAL 16
`define CVAL 17
`define MAXKVAL 9
`define TVPR 0.5
`define TRPR 0.5
